-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition"
-- CREATED		"Sat Feb 09 12:20:43 2019"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY SPIpulse1 IS 
	PORT
	(
		MISO :  IN  STD_LOGIC;
		CLK_50MHz :  IN  STD_LOGIC;
		CS :  OUT  STD_LOGIC;
		MSTR_CLK :  OUT  STD_LOGIC;
		MOSI :  OUT  STD_LOGIC
	);
END SPIpulse1;

ARCHITECTURE bdf_type OF SPIpulse1 IS 

COMPONENT spipulser
GENERIC (Count : INTEGER
			);
	PORT(CLK : IN STD_LOGIC;
		 input : IN STD_LOGIC;
		 output : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT addressblock
GENERIC (Count : INTEGER
			);
	PORT(CLK : IN STD_LOGIC;
		 NXTADD : IN STD_LOGIC;
		 ADDRESS : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT clk_divider
GENERIC (Count : INTEGER
			);
	PORT(CLK_IN : IN STD_LOGIC;
		 CLK_OUT : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT spi_master1
GENERIC (CPHA : STD_LOGIC;
			CPOL : STD_LOGIC;
			delay : INTEGER;
			dw : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 MISO : IN STD_LOGIC;
		 transmit : IN STD_LOGIC;
		 tx_data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 CS : OUT STD_LOGIC;
		 CLKO : OUT STD_LOGIC;
		 MOSI : OUT STD_LOGIC;
		 fPulse : OUT STD_LOGIC;
		 rx_data : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	CLK_1MHz :  STD_LOGIC;
SIGNAL	doneTx :  STD_LOGIC;
SIGNAL	pulseTx :  STD_LOGIC;
SIGNAL	rx :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(15 DOWNTO 0);


BEGIN 



b2v_inst : spipulser
GENERIC MAP(Count => 25
			)
PORT MAP(CLK => CLK_1MHz,
		 input => doneTx,
		 output => pulseTx);


b2v_inst2 : addressblock
GENERIC MAP(Count => 25
			)
PORT MAP(CLK => CLK_1MHz,
		 NXTADD => doneTx,
		 ADDRESS => SYNTHESIZED_WIRE_0);


b2v_inst20 : clk_divider
GENERIC MAP(Count => 25
			)
PORT MAP(CLK_IN => CLK_50MHz,
		 CLK_OUT => CLK_1MHz);


b2v_inst6 : spi_master1
GENERIC MAP(CPHA => '1',
			CPOL => '1',
			delay => 50,
			dw => 16
			)
PORT MAP(clk => CLK_1MHz,
		 MISO => MISO,
		 transmit => pulseTx,
		 tx_data => SYNTHESIZED_WIRE_0,
		 CS => CS,
		 CLKO => MSTR_CLK,
		 MOSI => MOSI,
		 fPulse => doneTx);


END bdf_type;